* minimal negative fixture placeholder
