* minimal borderline fixture placeholder
